`include "Lab5_Team1_Sliding_Window_Sequence_Detector.v"
`timescale 1ns / 1ps

module Sliding_Window_Sequence_Detector_t ();
    
endmodule