module test(in, out);
    input in;
    output out;
    not n1(out, in);
endmodule